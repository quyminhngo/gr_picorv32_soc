module PicoCounter (
    
);
endmodule